module cva6_tlb_DDFD6_A1F50 (
	clk_i,
	rst_ni,
	flush_i,
	flush_vvma_i,
	flush_gvma_i,
	s_st_enbl_i,
	g_st_enbl_i,
	v_i,
	update_i,
	lu_access_i,
	lu_asid_i,
	lu_vmid_i,
	lu_vaddr_i,
	lu_gpaddr_o,
	lu_content_o,
	lu_g_content_o,
	asid_to_be_flushed_i,
	vmid_to_be_flushed_i,
	vaddr_to_be_flushed_i,
	gpaddr_to_be_flushed_i,
	lu_is_page_o,
	lu_hit_o
);
	// removed localparam type pte_cva6_t_CVA6Cfg_type
	parameter [17102:0] pte_cva6_t_CVA6Cfg = 0;
	// removed localparam type tlb_update_cva6_t_CVA6Cfg_type
	// removed localparam type tlb_update_cva6_t_HYP_EXT_type
	// removed localparam type tlb_update_cva6_t_config_pkg_NrMaxRules_type
	parameter [17102:0] tlb_update_cva6_t_CVA6Cfg = 0;
	parameter [31:0] tlb_update_cva6_t_HYP_EXT = 0;
	parameter signed [31:0] tlb_update_cva6_t_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// Trace: core/cva6_mmu/cva6_tlb.sv:27:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/cva6_mmu/cva6_tlb.sv:28:20
	// removed localparam type pte_cva6_t
	// Trace: core/cva6_mmu/cva6_tlb.sv:29:20
	// removed localparam type tlb_update_cva6_t
	// Trace: core/cva6_mmu/cva6_tlb.sv:30:15
	parameter [31:0] TLB_ENTRIES = 4;
	// Trace: core/cva6_mmu/cva6_tlb.sv:31:15
	parameter [31:0] HYP_EXT = 0;
	// Trace: core/cva6_mmu/cva6_tlb.sv:33:5
	input wire clk_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:34:5
	input wire rst_ni;
	// Trace: core/cva6_mmu/cva6_tlb.sv:35:5
	input wire flush_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:36:5
	input wire flush_vvma_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:37:5
	input wire flush_gvma_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:38:5
	input wire s_st_enbl_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:39:5
	input wire g_st_enbl_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:40:5
	input wire v_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:42:5
	input wire [(((((((1 + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) >= ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) ? (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))))) + 1 : (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1)))) + 1)) + tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + ((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2))) + (((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9))) + (((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9))) - 1:0] update_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:44:5
	input wire lu_access_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:45:5
	input wire [CVA6Cfg[16940-:32] - 1:0] lu_asid_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:46:5
	input wire [CVA6Cfg[16908-:32] - 1:0] lu_vmid_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:47:5
	input wire [CVA6Cfg[17070-:32] - 1:0] lu_vaddr_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:48:5
	output reg [CVA6Cfg[17006-:32] - 1:0] lu_gpaddr_o;
	// Trace: core/cva6_mmu/cva6_tlb.sv:49:5
	output reg [(10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9:0] lu_content_o;
	// Trace: core/cva6_mmu/cva6_tlb.sv:50:5
	output reg [(10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9:0] lu_g_content_o;
	// Trace: core/cva6_mmu/cva6_tlb.sv:51:5
	input wire [CVA6Cfg[16940-:32] - 1:0] asid_to_be_flushed_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:52:5
	input wire [CVA6Cfg[16908-:32] - 1:0] vmid_to_be_flushed_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:53:5
	input wire [CVA6Cfg[17070-:32] - 1:0] vaddr_to_be_flushed_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:54:5
	input wire [CVA6Cfg[17006-:32] - 1:0] gpaddr_to_be_flushed_i;
	// Trace: core/cva6_mmu/cva6_tlb.sv:55:5
	output reg [CVA6Cfg[16011-:32] - 2:0] lu_is_page_o;
	// Trace: core/cva6_mmu/cva6_tlb.sv:56:5
	output reg lu_hit_o;
	// Trace: core/cva6_mmu/cva6_tlb.sv:58:3
	localparam GPPN2 = (CVA6Cfg[17102-:32] == 32 ? CVA6Cfg[17070-:32] - 33 : 10);
	// Trace: core/cva6_mmu/cva6_tlb.sv:60:3
	reg [((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (TLB_ENTRIES * (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1)) - 1 : (TLB_ENTRIES * (1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) - 1)):((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] tags_q;
	reg [((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (TLB_ENTRIES * (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1)) - 1 : (TLB_ENTRIES * (1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) - 1)):((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] tags_n;
	// Trace: core/cva6_mmu/cva6_tlb.sv:70:3
	reg [(TLB_ENTRIES * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) - 1:0] content_q;
	reg [(TLB_ENTRIES * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) - 1:0] content_n;
	// Trace: core/cva6_mmu/cva6_tlb.sv:76:3
	wire [(TLB_ENTRIES * CVA6Cfg[16011-:32]) - 1:0] vpn_match;
	// Trace: core/cva6_mmu/cva6_tlb.sv:77:3
	wire [(TLB_ENTRIES * CVA6Cfg[16011-:32]) - 1:0] level_match;
	// Trace: core/cva6_mmu/cva6_tlb.sv:78:3
	wire [((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? ((((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) - (HYP_EXT >= 0 ? 0 : HYP_EXT + 0)) + 1) * CVA6Cfg[16011-:32]) + (((HYP_EXT >= 0 ? 0 : HYP_EXT + 0) * CVA6Cfg[16011-:32]) - 1) : ((((HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1))) + 1) * CVA6Cfg[16011-:32]) + (((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) * CVA6Cfg[16011-:32]) - 1)):((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) * CVA6Cfg[16011-:32] : (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) * CVA6Cfg[16011-:32])] vaddr_vpn_match;
	// Trace: core/cva6_mmu/cva6_tlb.sv:79:3
	wire [((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? ((((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) - (HYP_EXT >= 0 ? 0 : HYP_EXT + 0)) + 1) * CVA6Cfg[16011-:32]) + (((HYP_EXT >= 0 ? 0 : HYP_EXT + 0) * CVA6Cfg[16011-:32]) - 1) : ((((HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1))) + 1) * CVA6Cfg[16011-:32]) + (((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) * CVA6Cfg[16011-:32]) - 1)):((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) * CVA6Cfg[16011-:32] : (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) * CVA6Cfg[16011-:32])] vaddr_level_match;
	// Trace: core/cva6_mmu/cva6_tlb.sv:80:3
	reg [TLB_ENTRIES - 1:0] lu_hit;
	// Trace: core/cva6_mmu/cva6_tlb.sv:81:3
	reg [TLB_ENTRIES - 1:0] replace_en;
	// Trace: core/cva6_mmu/cva6_tlb.sv:82:3
	reg [TLB_ENTRIES - 1:0] match_asid;
	// Trace: core/cva6_mmu/cva6_tlb.sv:83:3
	reg [TLB_ENTRIES - 1:0] match_vmid;
	// Trace: core/cva6_mmu/cva6_tlb.sv:84:3
	wire [(TLB_ENTRIES * CVA6Cfg[16011-:32]) - 1:0] page_match;
	// Trace: core/cva6_mmu/cva6_tlb.sv:85:3
	wire [((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? ((((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) - (HYP_EXT >= 0 ? 0 : HYP_EXT + 0)) + 1) * CVA6Cfg[16011-:32]) + (((HYP_EXT >= 0 ? 0 : HYP_EXT + 0) * CVA6Cfg[16011-:32]) - 1) : ((((HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1))) + 1) * CVA6Cfg[16011-:32]) + (((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) * CVA6Cfg[16011-:32]) - 1)):((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) * CVA6Cfg[16011-:32] : (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) * CVA6Cfg[16011-:32])] vpage_match;
	// Trace: core/cva6_mmu/cva6_tlb.sv:86:3
	wire [((CVA6Cfg[16011-:32] - 2) >= 0 ? (TLB_ENTRIES * (CVA6Cfg[16011-:32] - 1)) - 1 : (TLB_ENTRIES * (3 - CVA6Cfg[16011-:32])) + (CVA6Cfg[16011-:32] - 3)):((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2)] is_page_o;
	// Trace: core/cva6_mmu/cva6_tlb.sv:87:3
	reg [TLB_ENTRIES - 1:0] match_stage;
	// Trace: core/cva6_mmu/cva6_tlb.sv:88:3
	reg [(10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9:0] g_content;
	// Trace: core/cva6_mmu/cva6_tlb.sv:89:3
	reg [(TLB_ENTRIES * CVA6Cfg[387-:32]) - 1:0] gppn;
	// Trace: core/cva6_mmu/cva6_tlb.sv:90:3
	wire [2:0] v_st_enbl;
	// Trace: core/cva6_mmu/cva6_tlb.sv:92:3
	assign v_st_enbl = (CVA6Cfg[16543] ? {v_i, g_st_enbl_i, s_st_enbl_i} : {3 {1'sb1}});
	// Trace: core/cva6_mmu/cva6_tlb.sv:97:3
	genvar _gv_i_85;
	genvar _gv_x_2;
	genvar _gv_z_2;
	genvar _gv_w_2;
	// Trace: core/cva6_mmu/cva6_tlb.sv:98:3
	generate
		for (_gv_i_85 = 0; _gv_i_85 < TLB_ENTRIES; _gv_i_85 = _gv_i_85 + 1) begin : genblk1
			localparam i = _gv_i_85;
			for (_gv_x_2 = 0; _gv_x_2 < CVA6Cfg[16011-:32]; _gv_x_2 = _gv_x_2 + 1) begin : genblk1
				localparam x = _gv_x_2;
				// Trace: core/cva6_mmu/cva6_tlb.sv:102:9
				assign page_match[(i * CVA6Cfg[16011-:32]) + x] = (x == 0 ? 1 : ((HYP_EXT == 0) || (x == (CVA6Cfg[16011-:32] - 1)) ? &(tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)))) : (((((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT))))) - (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)))) : (((((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT))))) - (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + 1)) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)))) : (((((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT))))) - (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)))) : (((((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((HYP_EXT >= 0 ? 0 : HYP_EXT) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT))))) - (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + 1))) - (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + 1)+:(HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)] | ~v_st_enbl[HYP_EXT:0]) : (&v_st_enbl[HYP_EXT:0] ? (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))] && (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))))] || tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))))])) || (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))))] && (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 2) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 2) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))] || tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))])) : (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))] && s_st_enbl_i) || (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))))] && g_st_enbl_i))));
				// Trace: core/cva6_mmu/cva6_tlb.sv:110:9
				assign vpn_match[(i * CVA6Cfg[16011-:32]) + x] = ((CVA6Cfg[16543] && (x == (CVA6Cfg[16011-:32] - 1))) && ~s_st_enbl_i ? (lu_vaddr_i[(12 + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) * (x + 1))) - 1:12 + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) * x)] == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])))))) - (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + 1)+:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]]) && (lu_vaddr_i[12 + (HYP_EXT * (CVA6Cfg[16043-:32] - 1)):12 + (HYP_EXT * (CVA6Cfg[16043-:32] - (CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32])))] == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (((x + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? (CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT : (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + 1 : 1 - ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT))) - 1))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (((x + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? (CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT : (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + 1 : 1 - ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT))) - 1))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (((x + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? (CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT : (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + 1 : 1 - ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT))) - 1))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (((x + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? (CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT : (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + 1 : 1 - ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT))) - 1)))))) + (((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + 1 : 1 - ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT))) - 1)-:(((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) >= 0 ? ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT) + 1 : 1 - ((CVA6Cfg[16043-:32] % CVA6Cfg[16011-:32]) - HYP_EXT))]) : lu_vaddr_i[(12 + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) * (x + 1))) - 1:12 + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) * x)] == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])))))) - (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + 1)+:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]]);
				// Trace: core/cva6_mmu/cva6_tlb.sv:115:9
				assign level_match[(i * CVA6Cfg[16011-:32]) + x] = &vpn_match[(i * CVA6Cfg[16011-:32]) + ((CVA6Cfg[16011-:32] - 1) >= x ? CVA6Cfg[16011-:32] - 1 : ((CVA6Cfg[16011-:32] - 1) + ((CVA6Cfg[16011-:32] - 1) >= x ? ((CVA6Cfg[16011-:32] - 1) - x) + 1 : (x - (CVA6Cfg[16011-:32] - 1)) + 1)) - 1)-:((CVA6Cfg[16011-:32] - 1) >= x ? ((CVA6Cfg[16011-:32] - 1) - x) + 1 : (x - (CVA6Cfg[16011-:32] - 1)) + 1)] && page_match[(i * CVA6Cfg[16011-:32]) + x];
				for (_gv_z_2 = 0; _gv_z_2 < (HYP_EXT + 1); _gv_z_2 = _gv_z_2 + 1) begin : genblk1
					localparam z = _gv_z_2;
					// Trace: core/cva6_mmu/cva6_tlb.sv:119:11
					assign vpage_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + x] = (x == 0 ? 1 : tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (CVA6Cfg[16011-:32] - 1) - x : (CVA6Cfg[16011-:32] - 2) - ((CVA6Cfg[16011-:32] - 1) - x)) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z)))))]);
					// Trace: core/cva6_mmu/cva6_tlb.sv:120:11
					assign vaddr_level_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + x] = &vaddr_vpn_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + ((CVA6Cfg[16011-:32] - 1) >= x ? CVA6Cfg[16011-:32] - 1 : ((CVA6Cfg[16011-:32] - 1) + ((CVA6Cfg[16011-:32] - 1) >= x ? ((CVA6Cfg[16011-:32] - 1) - x) + 1 : (x - (CVA6Cfg[16011-:32] - 1)) + 1)) - 1)-:((CVA6Cfg[16011-:32] - 1) >= x ? ((CVA6Cfg[16011-:32] - 1) - x) + 1 : (x - (CVA6Cfg[16011-:32] - 1)) + 1)] && vpage_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? z : HYP_EXT - z)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + x];
				end
				// Trace: core/cva6_mmu/cva6_tlb.sv:124:9
				assign vaddr_vpn_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + x] = vaddr_to_be_flushed_i[(12 + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) * (x + 1))) - 1:12 + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) * x)] == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (x * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])))))) - (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + 1)+:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]];
			end
			if (CVA6Cfg[16543]) begin : genblk2
				// Trace: core/cva6_mmu/cva6_tlb.sv:132:9
				assign vaddr_vpn_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]] = gpaddr_to_be_flushed_i[20:12] == gppn[(i * CVA6Cfg[387-:32]) + 8-:9];
				// Trace: core/cva6_mmu/cva6_tlb.sv:133:9
				assign vaddr_vpn_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + HYP_EXT] = gpaddr_to_be_flushed_i[29:21] == gppn[(i * CVA6Cfg[387-:32]) + 17-:9];
				// Trace: core/cva6_mmu/cva6_tlb.sv:134:9
				assign vaddr_vpn_match[(((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]) + (HYP_EXT * 2)] = gpaddr_to_be_flushed_i[30 + GPPN2:30] == gppn[(i * CVA6Cfg[387-:32]) + ((18 + GPPN2) >= 18 ? 18 + GPPN2 : ((18 + GPPN2) + ((18 + GPPN2) >= 18 ? (18 + GPPN2) - 17 : 19 - (18 + GPPN2))) - 1)-:((18 + GPPN2) >= 18 ? (18 + GPPN2) - 17 : 19 - (18 + GPPN2))];
			end
			for (_gv_w_2 = 0; _gv_w_2 < (CVA6Cfg[16011-:32] - 1); _gv_w_2 = _gv_w_2 + 1) begin : genblk3
				localparam w = _gv_w_2;
				// Trace: core/cva6_mmu/cva6_tlb.sv:139:9
				assign is_page_o[(i * ((CVA6Cfg[16011-:32] - 2) >= 0 ? CVA6Cfg[16011-:32] - 1 : 3 - CVA6Cfg[16011-:32])) + ((CVA6Cfg[16011-:32] - 2) >= 0 ? w : (CVA6Cfg[16011-:32] - 2) - w)] = page_match[(i * CVA6Cfg[16011-:32]) + ((CVA6Cfg[16011-:32] - 1) - w)];
			end
		end
	endgenerate
	// Trace: core/cva6_mmu/cva6_tlb.sv:144:3
	function automatic [CVA6Cfg[17006-:32] - 1:0] sv2v_cast_8FFC6;
		input reg [CVA6Cfg[17006-:32] - 1:0] inp;
		sv2v_cast_8FFC6 = inp;
	endfunction
	function automatic [pte_cva6_t_CVA6Cfg[419-:32] - 1:0] sv2v_cast_5165A;
		input reg [pte_cva6_t_CVA6Cfg[419-:32] - 1:0] inp;
		sv2v_cast_5165A = inp;
	endfunction
	always @(*) begin : translation
		if (_sv2v_0)
			;
		// Trace: core/cva6_mmu/cva6_tlb.sv:147:5
		lu_hit = {TLB_ENTRIES {1'd0}};
		// Trace: core/cva6_mmu/cva6_tlb.sv:148:5
		lu_hit_o = 1'b0;
		// Trace: core/cva6_mmu/cva6_tlb.sv:149:5
		lu_content_o = {10'd0, sv2v_cast_5165A(0), 10'h000};
		// Trace: core/cva6_mmu/cva6_tlb.sv:150:5
		lu_g_content_o = {10'd0, sv2v_cast_5165A(0), 10'h000};
		// Trace: core/cva6_mmu/cva6_tlb.sv:151:5
		lu_is_page_o = {((CVA6Cfg[16011-:32] - 2) >= 0 ? CVA6Cfg[16011-:32] - 1 : 3 - CVA6Cfg[16011-:32]) {1'd0}};
		// Trace: core/cva6_mmu/cva6_tlb.sv:152:5
		match_asid = {TLB_ENTRIES {1'd0}};
		// Trace: core/cva6_mmu/cva6_tlb.sv:153:5
		match_vmid = (CVA6Cfg[16543] ? {TLB_ENTRIES {1'd0}} : {TLB_ENTRIES {1'd1}});
		// Trace: core/cva6_mmu/cva6_tlb.sv:154:5
		match_stage = {TLB_ENTRIES {1'd0}};
		// Trace: core/cva6_mmu/cva6_tlb.sv:155:5
		g_content = {10'd0, sv2v_cast_5165A(0), 10'h000};
		// Trace: core/cva6_mmu/cva6_tlb.sv:156:5
		lu_gpaddr_o = {CVA6Cfg[17006-:32] {1'd0}};
		// Trace: core/cva6_mmu/cva6_tlb.sv:158:5
		begin : sv2v_autoblock_1
			// Trace: core/cva6_mmu/cva6_tlb.sv:158:10
			reg [31:0] i;
			// Trace: core/cva6_mmu/cva6_tlb.sv:158:10
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin
					// Trace: core/cva6_mmu/cva6_tlb.sv:161:7
					match_asid[i] = (((lu_asid_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))))) + ((CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)) - 1)-:((CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg[16940-:32] + (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)]) || content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 4) : (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 5)]) && s_st_enbl_i) || !s_st_enbl_i;
					// Trace: core/cva6_mmu/cva6_tlb.sv:163:7
					if (CVA6Cfg[16543])
						// Trace: core/cva6_mmu/cva6_tlb.sv:164:9
						match_vmid[i] = ((lu_vmid_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg[16908-:32] + (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)]) && g_st_enbl_i) || !g_st_enbl_i;
					// Trace: core/cva6_mmu/cva6_tlb.sv:168:7
					match_stage[i] = tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) + (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1)) + 1 : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2))) + 1)) - 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) + (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1)) + 1 : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2))) + 1)) - 1)) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) + (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1)) + 1 : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2))) + 1)) - 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) + (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1)) + 1 : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2))) + 1)) - 1))) + (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1)) + 1 : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2))) + 1)) - 1)-:(((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) >= ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) ? (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1)) + 1 : (((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2))) + 1)] == v_st_enbl[HYP_EXT * 2:0];
					if (((tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] && match_asid[i]) && match_vmid[i]) && match_stage[i]) begin
						// Trace: core/cva6_mmu/cva6_tlb.sv:172:9
						if (CVA6Cfg[16543] && vpn_match[(i * CVA6Cfg[16011-:32]) + (HYP_EXT * 2)]) begin
							begin
								// Trace: core/cva6_mmu/cva6_tlb.sv:173:11
								if (s_st_enbl_i) begin
									// Trace: core/cva6_mmu/cva6_tlb.sv:174:13
									lu_gpaddr_o = {content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) >= (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) ? (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) >= (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1 : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1)) - 1)-:((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) >= (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1 : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1)], lu_vaddr_i[11:0]};
									// Trace: core/cva6_mmu/cva6_tlb.sv:176:13
									if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))])
										// Trace: core/cva6_mmu/cva6_tlb.sv:177:15
										lu_gpaddr_o[(12 + ((2 * CVA6Cfg[16043-:32]) / CVA6Cfg[16011-:32])) - 1:12] = lu_vaddr_i[(12 + ((2 * CVA6Cfg[16043-:32]) / CVA6Cfg[16011-:32])) - 1:12];
									if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))])
										// Trace: core/cva6_mmu/cva6_tlb.sv:180:15
										lu_gpaddr_o[(12 + (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1:12] = lu_vaddr_i[(12 + (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1:12];
								end
								else
									// Trace: core/cva6_mmu/cva6_tlb.sv:182:13
									lu_gpaddr_o = sv2v_cast_8FFC6(lu_vaddr_i[(CVA6Cfg[17102-:32] == 32 ? CVA6Cfg[17070-:32] : CVA6Cfg[17006-:32]) - 1:0]);
							end
						end
						if (|level_match[i * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]]) begin
							// Trace: core/cva6_mmu/cva6_tlb.sv:187:11
							lu_is_page_o = is_page_o[((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) + (i * ((CVA6Cfg[16011-:32] - 2) >= 0 ? CVA6Cfg[16011-:32] - 1 : 3 - CVA6Cfg[16011-:32]))+:((CVA6Cfg[16011-:32] - 2) >= 0 ? CVA6Cfg[16011-:32] - 1 : 3 - CVA6Cfg[16011-:32])];
							// Trace: core/cva6_mmu/cva6_tlb.sv:188:11
							lu_content_o = content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))-:(((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) >= ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) ? (((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)) + 1 : (((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) - ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))) + 1)];
							// Trace: core/cva6_mmu/cva6_tlb.sv:189:11
							lu_hit_o = 1'b1;
							// Trace: core/cva6_mmu/cva6_tlb.sv:190:11
							lu_hit[i] = 1'b1;
							// Trace: core/cva6_mmu/cva6_tlb.sv:192:11
							if (CVA6Cfg[16543]) begin
								// Trace: core/cva6_mmu/cva6_tlb.sv:194:13
								g_content = content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)-:(((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9))];
								// Trace: core/cva6_mmu/cva6_tlb.sv:195:13
								if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))))])
									// Trace: core/cva6_mmu/cva6_tlb.sv:195:54
									g_content[(pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 9):(pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1)] = lu_gpaddr_o[20:12];
								if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)))))])
									// Trace: core/cva6_mmu/cva6_tlb.sv:196:48
									g_content[(pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 18):(pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1)] = lu_gpaddr_o[29:12];
								// Trace: core/cva6_mmu/cva6_tlb.sv:198:13
								lu_g_content_o = (level_match[(i * CVA6Cfg[16011-:32]) + (CVA6Cfg[16011-:32] - 1)] ? content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)-:(((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9))] : g_content);
							end
						end
					end
				end
		end
	end
	// Trace: core/cva6_mmu/cva6_tlb.sv:205:3
	wire [HYP_EXT:0] asid_to_be_flushed_is0;
	// Trace: core/cva6_mmu/cva6_tlb.sv:206:3
	wire [HYP_EXT:0] vaddr_to_be_flushed_is0;
	// Trace: core/cva6_mmu/cva6_tlb.sv:207:3
	wire vmid_to_be_flushed_is0;
	// Trace: core/cva6_mmu/cva6_tlb.sv:208:3
	wire gpaddr_to_be_flushed_is0;
	// Trace: core/cva6_mmu/cva6_tlb.sv:210:3
	assign asid_to_be_flushed_is0 = ~(|asid_to_be_flushed_i);
	// Trace: core/cva6_mmu/cva6_tlb.sv:211:3
	assign vaddr_to_be_flushed_is0 = ~(|vaddr_to_be_flushed_i);
	// Trace: core/cva6_mmu/cva6_tlb.sv:212:3
	assign vmid_to_be_flushed_is0 = ~(|vmid_to_be_flushed_i);
	// Trace: core/cva6_mmu/cva6_tlb.sv:213:3
	assign gpaddr_to_be_flushed_is0 = ~(|gpaddr_to_be_flushed_i);
	// Trace: core/cva6_mmu/cva6_tlb.sv:218:3
	function automatic [CVA6Cfg[16043-:32] - 1:0] sv2v_cast_4DD5A;
		input reg [CVA6Cfg[16043-:32] - 1:0] inp;
		sv2v_cast_4DD5A = inp;
	endfunction
	function automatic [((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1:0] sv2v_cast_77756;
		input reg [((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1:0] inp;
		sv2v_cast_77756 = inp;
	endfunction
	always @(*) begin : update_flush
		if (_sv2v_0)
			;
		// Trace: core/cva6_mmu/cva6_tlb.sv:219:5
		tags_n = tags_q;
		// Trace: core/cva6_mmu/cva6_tlb.sv:220:5
		content_n = content_q;
		// Trace: core/cva6_mmu/cva6_tlb.sv:222:5
		begin : sv2v_autoblock_2
			// Trace: core/cva6_mmu/cva6_tlb.sv:222:10
			reg [31:0] i;
			// Trace: core/cva6_mmu/cva6_tlb.sv:222:10
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin
					// Trace: core/cva6_mmu/cva6_tlb.sv:225:7
					if (CVA6Cfg[16543]) begin
						begin
							// Trace: core/cva6_mmu/cva6_tlb.sv:227:9
							if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1))]) begin
								// Trace: core/cva6_mmu/cva6_tlb.sv:228:11
								gppn[i * CVA6Cfg[387-:32]+:CVA6Cfg[387-:32]] = content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) >= (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) ? (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) >= (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1 : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1)) - 1)-:((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) >= (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1 : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - (pte_cva6_t_CVA6Cfg[419-:32] - 1))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (pte_cva6_t_CVA6Cfg[419-:32] + 9))) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] + 9) - ((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)))) : ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) + (((pte_cva6_t_CVA6Cfg[419-:32] - 1) - (CVA6Cfg[387-:32] - 1)) - (pte_cva6_t_CVA6Cfg[419-:32] + 9)))) + 1)];
								// Trace: core/cva6_mmu/cva6_tlb.sv:229:11
								if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? HYP_EXT : (CVA6Cfg[16011-:32] - 2) - HYP_EXT) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))])
									// Trace: core/cva6_mmu/cva6_tlb.sv:230:13
									gppn[(i * CVA6Cfg[387-:32]) + ((CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]) - 1)-:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]] = tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1)))) - (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + 1)+:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]];
								if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) - (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT))) : (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? 0 : CVA6Cfg[16011-:32] - 2) * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)))))])
									// Trace: core/cva6_mmu/cva6_tlb.sv:232:13
									gppn[(i * CVA6Cfg[387-:32]) + ((2 * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1)-:2 * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])] = {tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (HYP_EXT * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (HYP_EXT * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (HYP_EXT * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) - (HYP_EXT * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])))))) - (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + 1)+:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]], tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) - 1)))) - (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + 1)+:CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]]};
							end
							else
								// Trace: core/cva6_mmu/cva6_tlb.sv:236:11
								gppn[(i * CVA6Cfg[387-:32]) + (CVA6Cfg[16043-:32] - 1)-:CVA6Cfg[16043-:32]] = sv2v_cast_4DD5A(tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) >= ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)) ? ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) + 1 : (((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) + 1)) - 1)-:((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) >= ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)) ? ((((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) - ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) + 1 : (((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)) - (((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32])) + ((((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) + 1)]);
						end
					end
					if (flush_i) begin
						begin
							// Trace: core/cva6_mmu/cva6_tlb.sv:242:9
							if (!tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)))] || (HYP_EXT == 0)) begin
								begin
									// Trace: core/cva6_mmu/cva6_tlb.sv:245:11
									if (asid_to_be_flushed_is0 && vaddr_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:245:66
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if ((asid_to_be_flushed_is0 && |vaddr_level_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]]) && ~vaddr_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:248:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if ((((!content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 4) : (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 5)] && |vaddr_level_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]]) && (asid_to_be_flushed_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))))) + ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)) - 1)-:((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)])) && !vaddr_to_be_flushed_is0) && !asid_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:251:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if (((!content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 4) : (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 5)] && vaddr_to_be_flushed_is0) && (asid_to_be_flushed_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))))) + ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)) - 1)-:((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)])) && !asid_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:254:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
								end
							end
						end
					end
					else if (flush_vvma_i && CVA6Cfg[16543]) begin
						begin
							// Trace: core/cva6_mmu/cva6_tlb.sv:257:9
							if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - (HYP_EXT * 2)) : 1 - (HYP_EXT * 2)))] && tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - (HYP_EXT * 2) : 1))]) begin
								begin
									// Trace: core/cva6_mmu/cva6_tlb.sv:260:11
									if ((asid_to_be_flushed_is0 && vaddr_to_be_flushed_is0) && ((tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))] && (lu_vmid_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)])) || !tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))]))
										// Trace: core/cva6_mmu/cva6_tlb.sv:261:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if (((asid_to_be_flushed_is0 && |vaddr_level_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]]) && ~vaddr_to_be_flushed_is0) && ((tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))] && (lu_vmid_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)])) || !tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))]))
										// Trace: core/cva6_mmu/cva6_tlb.sv:264:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if ((((!content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 4) : (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 5)] && |vaddr_level_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? 0 : HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]]) && ((asid_to_be_flushed_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))))) + ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)) - 1)-:((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)]) && ((tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))] && (lu_vmid_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)])) || !tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))]))) && !vaddr_to_be_flushed_is0) && !asid_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:267:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if (((!content_q[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 4) : (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 5)] && vaddr_to_be_flushed_is0) && ((asid_to_be_flushed_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))))) + ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)) - 1)-:((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) >= (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) ? ((CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))))) + 1 : ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) - (CVA6Cfg.ASID_WIDTH + (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + 1)]) && ((tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))] && (lu_vmid_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)])) || !tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))]))) && !asid_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:270:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
								end
							end
						end
					end
					else if (flush_gvma_i && CVA6Cfg[16543]) begin
						begin
							// Trace: core/cva6_mmu/cva6_tlb.sv:273:9
							if (tags_q[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - ((HYP_EXT * 2) >= 0 ? (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0) - ((HYP_EXT * 2) - HYP_EXT) : 1 - HYP_EXT))]) begin
								begin
									// Trace: core/cva6_mmu/cva6_tlb.sv:276:11
									if (vmid_to_be_flushed_is0 && gpaddr_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:276:67
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if ((vmid_to_be_flushed_is0 && |vaddr_level_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]]) && ~gpaddr_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:279:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if (((|vaddr_level_match[((HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)) >= (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) ? (i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT) : (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) - (((i * (HYP_EXT >= 0 ? HYP_EXT + 1 : 1 - HYP_EXT)) + (HYP_EXT >= 0 ? HYP_EXT : HYP_EXT - HYP_EXT)) - (HYP_EXT >= 0 ? (TLB_ENTRIES * (HYP_EXT + 1)) - 1 : (TLB_ENTRIES * (1 - HYP_EXT)) + (HYP_EXT - 1)))) * CVA6Cfg[16011-:32]+:CVA6Cfg[16011-:32]] && (vmid_to_be_flushed_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)])) && ~gpaddr_to_be_flushed_is0) && ~vmid_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:282:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
									else if ((gpaddr_to_be_flushed_is0 && (vmid_to_be_flushed_i == tags_q[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) : (((i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))) : (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))))) + ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)) - 1)-:((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) >= (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) ? ((CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0)))) - (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1)))) + 1 : ((((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 1))) - (CVA6Cfg.VMID_WIDTH + (((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels)) + ((((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1) + (((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2)) + 0))))) + 1)])) && !vmid_to_be_flushed_is0)
										// Trace: core/cva6_mmu/cva6_tlb.sv:285:13
										tags_n[(i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))) + ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)] = 1'b0;
								end
							end
						end
					end
					else if ((update_i[1 + ((((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) >= ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) ? (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))))) + 1 : (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1)))) + 1) + (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))))))] & replace_en[i]) & !lu_hit_o) begin
						// Trace: core/cva6_mmu/cva6_tlb.sv:290:9
						tags_n[((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? 0 : ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) + (i * ((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)))+:((((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg[16940-:32] + CVA6Cfg[16908-:32]) + ((CVA6Cfg[16011-:32] + HYP_EXT) * (CVA6Cfg[16043-:32] / CVA6Cfg[16011-:32]))) + (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg[16011-:32] - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg[16011-:32] - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg[16011-:32] - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg[16011-:32]) * (HYP_EXT + 1)) + (((CVA6Cfg[16011-:32] - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg[16011-:32]) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg[16011-:32] - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0))] = {update_i[tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))-:((tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))) >= (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)))) ? ((tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))) - (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))))) + 1 : ((tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)))) - (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))))) + 1)], update_i[tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))-:((tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))) >= (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))) ? ((tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))) - (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)))) + 1 : ((((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))) - (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))) + 1)], sv2v_cast_77756(update_i[tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))))-:((tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))))) >= (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))))) ? ((tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))))) - (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)))))) + 1 : ((tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))))) - (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))))) + 1)]), update_i[(((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) >= ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) ? (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))))) + 1 : (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1)))) + 1) + (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))))-:(((((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) >= ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) ? (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))))) + 1 : (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1)))) + 1) + (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))))) >= (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)))))) ? (((((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) >= ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) ? (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))))) + 1 : (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1)))) + 1) + (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))))))) - (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))))))) + 1 : ((tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)))))) - ((((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) >= ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) ? (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))))) + 1 : (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? 0 : tlb_update_cva6_t_HYP_EXT + 0) : (tlb_update_cva6_t_HYP_EXT >= 0 ? (tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1) : tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT)))) - ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT >= 0 ? ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1 : ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) * (1 - tlb_update_cva6_t_HYP_EXT)) + (tlb_update_cva6_t_HYP_EXT - 1)) : (tlb_update_cva6_t_HYP_EXT >= 0 ? ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (tlb_update_cva6_t_HYP_EXT + 1)) + (((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (tlb_update_cva6_t_HYP_EXT + 1)) - 1) : ((3 - tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (1 - tlb_update_cva6_t_HYP_EXT)) + ((tlb_update_cva6_t_HYP_EXT + ((tlb_update_cva6_t_CVA6Cfg[8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8418 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2) * (1 - tlb_update_cva6_t_HYP_EXT))) - 1)))) + 1) + (tlb_update_cva6_t_CVA6Cfg[8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8450 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8482 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9379 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (tlb_update_cva6_t_CVA6Cfg[9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9315 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9347 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + (32 + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + ((tlb_update_cva6_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))))))) + 1)], update_i[((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))-:((((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))) >= ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)) ? ((((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))) - ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0))) + 1 : (((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)) - (((tlb_update_cva6_t_HYP_EXT * 2) >= 0 ? (tlb_update_cva6_t_HYP_EXT * 2) + 1 : 1 - (tlb_update_cva6_t_HYP_EXT * 2)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)))) + 1)], 1'b1};
						// Trace: core/cva6_mmu/cva6_tlb.sv:299:9
						content_n[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))-:(((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) >= ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) ? (((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)) + 1 : (((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) - ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))) + 1)] = update_i[(((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)-:(((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) >= ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) ? (((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)) - ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0)) + 1 : (((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + 0) - ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) + ((((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1))) + 1)];
						// Trace: core/cva6_mmu/cva6_tlb.sv:300:9
						if (CVA6Cfg[16543])
							// Trace: core/cva6_mmu/cva6_tlb.sv:300:26
							content_n[(i * ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)))) + ((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1)-:(((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9))] = update_i[(((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9)) - 1-:(((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + tlb_update_cva6_t_CVA6Cfg[419-:32]) + 9))];
					end
				end
		end
	end
	// Trace: core/cva6_mmu/cva6_tlb.sv:308:3
	reg [(2 * (TLB_ENTRIES - 1)) - 1:0] plru_tree_q;
	reg [(2 * (TLB_ENTRIES - 1)) - 1:0] plru_tree_n;
	// Trace: core/cva6_mmu/cva6_tlb.sv:309:3
	always @(*) begin : plru_replacement
		if (_sv2v_0)
			;
		// Trace: core/cva6_mmu/cva6_tlb.sv:310:5
		plru_tree_n = plru_tree_q;
		// Trace: core/cva6_mmu/cva6_tlb.sv:334:1
		begin : sv2v_autoblock_3
			// Trace: core/cva6_mmu/cva6_tlb.sv:335:9
			reg [31:0] i;
			// Trace: core/cva6_mmu/cva6_tlb.sv:335:9
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin : sv2v_autoblock_4
					// Trace: core/cva6_mmu/cva6_tlb.sv:337:7
					reg [31:0] idx_base;
					reg [31:0] shift;
					reg [31:0] new_index;
					// Trace: core/cva6_mmu/cva6_tlb.sv:339:7
					if (lu_hit[i] & lu_access_i)
						// Trace: core/cva6_mmu/cva6_tlb.sv:341:9
						begin : sv2v_autoblock_5
							// Trace: core/cva6_mmu/cva6_tlb.sv:341:14
							reg [31:0] lvl;
							// Trace: core/cva6_mmu/cva6_tlb.sv:341:14
							for (lvl = 0; lvl < $clog2(TLB_ENTRIES); lvl = lvl + 1)
								begin
									// Trace: core/cva6_mmu/cva6_tlb.sv:342:11
									idx_base = $unsigned((2 ** lvl) - 1);
									// Trace: core/cva6_mmu/cva6_tlb.sv:344:11
									shift = $clog2(TLB_ENTRIES) - lvl;
									// Trace: core/cva6_mmu/cva6_tlb.sv:346:11
									new_index = ~((i >> (shift - 1)) & 32'b00000000000000000000000000000001);
									// Trace: core/cva6_mmu/cva6_tlb.sv:347:11
									plru_tree_n[idx_base + (i >> shift)] = new_index[0];
								end
						end
				end
		end
		begin : sv2v_autoblock_6
			// Trace: core/cva6_mmu/cva6_tlb.sv:365:10
			reg [31:0] i;
			// Trace: core/cva6_mmu/cva6_tlb.sv:365:10
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin : sv2v_autoblock_7
					// Trace: core/cva6_mmu/cva6_tlb.sv:366:7
					reg en;
					// Trace: core/cva6_mmu/cva6_tlb.sv:367:7
					reg [31:0] idx_base;
					reg [31:0] shift;
					reg [31:0] new_index;
					// Trace: core/cva6_mmu/cva6_tlb.sv:368:7
					en = 1'b1;
					// Trace: core/cva6_mmu/cva6_tlb.sv:369:7
					begin : sv2v_autoblock_8
						// Trace: core/cva6_mmu/cva6_tlb.sv:369:12
						reg [31:0] lvl;
						// Trace: core/cva6_mmu/cva6_tlb.sv:369:12
						for (lvl = 0; lvl < $clog2(TLB_ENTRIES); lvl = lvl + 1)
							begin
								// Trace: core/cva6_mmu/cva6_tlb.sv:370:9
								idx_base = $unsigned((2 ** lvl) - 1);
								// Trace: core/cva6_mmu/cva6_tlb.sv:372:9
								shift = $clog2(TLB_ENTRIES) - lvl;
								// Trace: core/cva6_mmu/cva6_tlb.sv:375:9
								new_index = (i >> (shift - 1)) & 32'b00000000000000000000000000000001;
								// Trace: core/cva6_mmu/cva6_tlb.sv:376:9
								if (new_index[0])
									// Trace: core/cva6_mmu/cva6_tlb.sv:377:11
									en = en & plru_tree_q[idx_base + (i >> shift)];
								else
									// Trace: core/cva6_mmu/cva6_tlb.sv:379:11
									en = en & ~plru_tree_q[idx_base + (i >> shift)];
							end
					end
					// Trace: core/cva6_mmu/cva6_tlb.sv:382:7
					replace_en[i] = en;
				end
		end
	end
	// Trace: core/cva6_mmu/cva6_tlb.sv:387:3
	function automatic [((((((CVA6Cfg.ASID_WIDTH + CVA6Cfg.VMID_WIDTH) + ((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels))) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg.ASID_WIDTH + CVA6Cfg.VMID_WIDTH) + ((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels))) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg.ASID_WIDTH + CVA6Cfg.VMID_WIDTH) + ((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels))) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)) - 1:0] sv2v_cast_27262;
		input reg [((((((CVA6Cfg.ASID_WIDTH + CVA6Cfg.VMID_WIDTH) + ((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels))) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0) >= 0 ? ((((CVA6Cfg.ASID_WIDTH + CVA6Cfg.VMID_WIDTH) + ((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels))) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 1 : 1 - (((((CVA6Cfg.ASID_WIDTH + CVA6Cfg.VMID_WIDTH) + ((CVA6Cfg.PtLevels + HYP_EXT) * (CVA6Cfg.VpnLen / CVA6Cfg.PtLevels))) + (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) >= ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) ? (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))))) + 1 : (((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? 0 : HYP_EXT + 0) : (HYP_EXT >= 0 ? (CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1) : HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT)))) - ((CVA6Cfg.PtLevels - 2) >= 0 ? (HYP_EXT >= 0 ? ((CVA6Cfg.PtLevels - 1) * (HYP_EXT + 1)) - 1 : ((CVA6Cfg.PtLevels - 1) * (1 - HYP_EXT)) + (HYP_EXT - 1)) : (HYP_EXT >= 0 ? ((3 - CVA6Cfg.PtLevels) * (HYP_EXT + 1)) + (((CVA6Cfg.PtLevels - 2) * (HYP_EXT + 1)) - 1) : ((3 - CVA6Cfg.PtLevels) * (1 - HYP_EXT)) + ((HYP_EXT + ((CVA6Cfg.PtLevels - 2) * (1 - HYP_EXT))) - 1)))) + 1)) + ((HYP_EXT * 2) >= 0 ? (HYP_EXT * 2) + 1 : 1 - (HYP_EXT * 2))) + 0)) - 1:0] inp;
		sv2v_cast_27262 = inp;
	endfunction
	function automatic [((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9))) - 1:0] sv2v_cast_6265D;
		input reg [((((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9)) + (((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9) >= 0 ? (10 + pte_cva6_t_CVA6Cfg[419-:32]) + 10 : 1 - ((10 + pte_cva6_t_CVA6Cfg[419-:32]) + 9))) - 1:0] inp;
		sv2v_cast_6265D = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni)
		// Trace: core/cva6_mmu/cva6_tlb.sv:388:5
		if (~rst_ni) begin
			// Trace: core/cva6_mmu/cva6_tlb.sv:389:7
			tags_q <= {TLB_ENTRIES {sv2v_cast_27262(0)}};
			// Trace: core/cva6_mmu/cva6_tlb.sv:390:7
			content_q <= {TLB_ENTRIES {sv2v_cast_6265D(0)}};
			// Trace: core/cva6_mmu/cva6_tlb.sv:391:7
			plru_tree_q <= {2 * (TLB_ENTRIES - 1) {1'd0}};
		end
		else begin
			// Trace: core/cva6_mmu/cva6_tlb.sv:393:7
			tags_q <= tags_n;
			// Trace: core/cva6_mmu/cva6_tlb.sv:394:7
			content_q <= content_n;
			// Trace: core/cva6_mmu/cva6_tlb.sv:395:7
			plru_tree_q <= plru_tree_n;
		end
	// Trace: core/cva6_mmu/cva6_tlb.sv:405:3
	initial begin : p_assertions
		// Trace: core/cva6_mmu/cva6_tlb.sv:406:5
	end
	// Trace: core/cva6_mmu/cva6_tlb.sv:419:3
	function signed [31:0] countSetBits;
		// Trace: core/cva6_mmu/cva6_tlb.sv:419:29
		input reg [TLB_ENTRIES - 1:0] vector;
		// Trace: core/cva6_mmu/cva6_tlb.sv:420:5
		reg signed [31:0] count;
		begin
			count = 0;
			// Trace: core/cva6_mmu/cva6_tlb.sv:421:5
			begin : sv2v_autoblock_9
				integer idx;
				for (idx = TLB_ENTRIES - 1; idx >= 0; idx = idx - 1)
					begin
						// Trace: core/cva6_mmu/cva6_tlb.sv:422:7
						count = count + vector[idx];
					end
			end
			countSetBits = count;
		end
	endfunction
	// Trace: core/cva6_mmu/cva6_tlb.sv:427:3
	// removed an assertion item
	// assert property (@(posedge clk_i) 
	// 	countSetBits(lu_hit) <= 1
	// ) else begin
	// 	// Trace: core/cva6_mmu/cva6_tlb.sv:429:5
	// 	$error("More then one hit in TLB!");
	// 	// Trace: core/cva6_mmu/cva6_tlb.sv:430:5
	// 	$stop;
	// end
	// Trace: core/cva6_mmu/cva6_tlb.sv:432:3
	// removed an assertion item
	// assert property (@(posedge clk_i) 
	// 	countSetBits(replace_en) <= 1
	// ) else begin
	// 	// Trace: core/cva6_mmu/cva6_tlb.sv:434:5
	// 	$error("More then one TLB entry selected for next replace!");
	// 	// Trace: core/cva6_mmu/cva6_tlb.sv:435:5
	// 	$stop;
	// end
	initial _sv2v_0 = 0;
endmodule
