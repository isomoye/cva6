module unread (d_i);
	// Trace: vendor/pulp-platform/common_cells/src/unread.sv:17:5
	input wire d_i;
endmodule
